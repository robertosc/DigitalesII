`timescale 	1ns	/ 100ps
`include "alarma_desc_conductual.v"

module Pruebas; 
	alarma_desc_conductual	cond(/*AUTOINST*/);
   
endmodule
